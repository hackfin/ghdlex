vfx2fifo.vhdl